module cpu (

);

endmodule